VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_2kbyte_1rw1r_32x512_8
   CLASS BLOCK ;
   FOREIGN sky130_sram_2kbyte_1rw1r_32x512_8 ;
   SIZE 683.1 BY 416.54 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.04 0.0 121.42 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.6 0.0 132.98 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 0.0 190.78 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 0.0 214.58 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 0.0 256.06 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  85.68 0.0 86.06 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.76 1.06 141.14 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 1.06 149.98 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.04 1.06 155.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.88 1.06 164.26 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 1.06 169.02 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 179.52 1.06 179.9 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.28 1.06 184.66 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  598.4 415.48 598.78 416.54 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  592.28 415.48 592.66 416.54 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 96.56 683.1 96.94 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 88.4 683.1 88.78 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 81.6 683.1 81.98 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 74.12 683.1 74.5 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 68.0 683.1 68.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.08 0.0 616.46 1.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.76 0.0 617.14 1.06 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 1.06 40.5 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 395.76 683.1 396.14 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 49.64 1.06 50.02 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 41.48 1.06 41.86 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  654.16 415.48 654.54 416.54 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.12 0.0 91.5 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.92 0.0 98.3 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.68 0.0 103.06 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.8 0.0 109.18 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 0.0 168.34 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 0.0 268.3 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 0.0 280.54 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 0.0 317.94 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.8 0.0 330.18 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 0.0 355.34 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 0.0 367.58 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 0.0 379.82 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  392.36 0.0 392.74 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 0.0 417.9 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 0.0 430.14 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.68 0.0 443.06 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 0.0 455.3 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.16 0.0 467.54 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  479.4 0.0 479.78 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 0.0 492.7 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  504.56 0.0 504.94 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 0.0 517.18 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  529.72 0.0 530.1 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 415.48 143.86 416.54 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 415.48 155.42 416.54 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 415.48 167.66 416.54 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 415.48 181.26 416.54 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 415.48 192.82 416.54 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 415.48 205.74 416.54 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 415.48 217.98 416.54 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 415.48 230.9 416.54 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 415.48 243.14 416.54 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 415.48 256.06 416.54 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 415.48 268.3 416.54 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 415.48 281.22 416.54 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 415.48 292.78 416.54 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 415.48 305.02 416.54 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.24 415.48 318.62 416.54 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 415.48 330.86 416.54 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 415.48 343.1 416.54 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 415.48 355.34 416.54 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 415.48 368.26 416.54 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 415.48 379.82 416.54 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 415.48 393.42 416.54 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 415.48 405.66 416.54 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 415.48 417.9 416.54 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 415.48 430.14 416.54 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 415.48 442.38 416.54 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 415.48 455.3 416.54 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.84 415.48 468.22 416.54 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.08 415.48 480.46 416.54 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 415.48 492.7 416.54 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 415.48 505.62 416.54 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 415.48 517.18 416.54 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.4 415.48 530.78 416.54 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 411.78 ;
         LAYER met4 ;
         RECT  676.6 4.76 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 410.04 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 4.76 678.34 6.5 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  680.0 1.36 681.74 415.18 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 415.18 ;
         LAYER met3 ;
         RECT  1.36 1.36 681.74 3.1 ;
         LAYER met3 ;
         RECT  1.36 413.44 681.74 415.18 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met2 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met3 ;
      RECT  1.66 140.16 682.48 141.74 ;
      RECT  0.62 141.74 1.66 149.0 ;
      RECT  0.62 150.58 1.66 154.44 ;
      RECT  0.62 156.02 1.66 163.28 ;
      RECT  0.62 164.86 1.66 168.04 ;
      RECT  0.62 169.62 1.66 178.92 ;
      RECT  0.62 180.5 1.66 183.68 ;
      RECT  1.66 95.96 681.44 97.54 ;
      RECT  1.66 97.54 681.44 140.16 ;
      RECT  681.44 97.54 682.48 140.16 ;
      RECT  681.44 89.38 682.48 95.96 ;
      RECT  681.44 82.58 682.48 87.8 ;
      RECT  681.44 75.1 682.48 81.0 ;
      RECT  681.44 68.98 682.48 73.52 ;
      RECT  1.66 141.74 681.44 395.16 ;
      RECT  1.66 395.16 681.44 396.74 ;
      RECT  681.44 141.74 682.48 395.16 ;
      RECT  0.62 50.62 1.66 140.16 ;
      RECT  0.62 42.46 1.66 49.04 ;
      RECT  1.66 396.74 4.16 409.44 ;
      RECT  1.66 409.44 4.16 412.38 ;
      RECT  4.16 396.74 678.94 409.44 ;
      RECT  678.94 396.74 681.44 409.44 ;
      RECT  678.94 409.44 681.44 412.38 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 95.96 ;
      RECT  4.16 7.1 678.94 95.96 ;
      RECT  678.94 4.16 681.44 7.1 ;
      RECT  678.94 7.1 681.44 95.96 ;
      RECT  681.44 0.62 682.34 0.76 ;
      RECT  681.44 3.7 682.34 67.4 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 3.7 ;
      RECT  682.34 3.7 682.48 67.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 39.52 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 39.52 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 678.94 0.76 ;
      RECT  4.16 3.7 678.94 4.16 ;
      RECT  678.94 0.62 681.44 0.76 ;
      RECT  678.94 3.7 681.44 4.16 ;
      RECT  0.62 185.26 0.76 412.84 ;
      RECT  0.62 412.84 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 185.26 1.66 412.84 ;
      RECT  0.76 415.78 1.66 415.92 ;
      RECT  681.44 396.74 682.34 412.84 ;
      RECT  681.44 415.78 682.34 415.92 ;
      RECT  682.34 396.74 682.48 412.84 ;
      RECT  682.34 412.84 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  1.66 412.38 4.16 412.84 ;
      RECT  1.66 415.78 4.16 415.92 ;
      RECT  4.16 412.38 678.94 412.84 ;
      RECT  4.16 415.78 678.94 415.92 ;
      RECT  678.94 412.38 681.44 412.84 ;
      RECT  678.94 415.78 681.44 415.92 ;
   LAYER  met4 ;
      RECT  115.0 1.66 116.58 415.92 ;
      RECT  116.58 0.62 120.44 1.66 ;
      RECT  122.02 0.62 126.56 1.66 ;
      RECT  128.14 0.62 132.0 1.66 ;
      RECT  133.58 0.62 137.44 1.66 ;
      RECT  144.46 0.62 149.68 1.66 ;
      RECT  157.38 0.62 161.24 1.66 ;
      RECT  162.82 0.62 166.68 1.66 ;
      RECT  173.7 0.62 178.92 1.66 ;
      RECT  185.94 0.62 189.8 1.66 ;
      RECT  198.18 0.62 202.72 1.66 ;
      RECT  209.74 0.62 213.6 1.66 ;
      RECT  220.62 0.62 225.84 1.66 ;
      RECT  232.86 0.62 237.4 1.66 ;
      RECT  244.42 0.62 248.28 1.66 ;
      RECT  256.66 0.62 260.52 1.66 ;
      RECT  262.1 0.62 265.96 1.66 ;
      RECT  272.98 0.62 278.2 1.66 ;
      RECT  285.9 0.62 289.76 1.66 ;
      RECT  81.22 0.62 85.08 1.66 ;
      RECT  116.58 1.66 597.8 414.88 ;
      RECT  597.8 1.66 599.38 414.88 ;
      RECT  593.26 414.88 597.8 415.92 ;
      RECT  599.38 414.88 653.56 415.92 ;
      RECT  86.66 0.62 90.52 1.66 ;
      RECT  92.1 0.62 97.32 1.66 ;
      RECT  98.9 0.62 102.08 1.66 ;
      RECT  103.66 0.62 108.2 1.66 ;
      RECT  109.78 0.62 115.0 1.66 ;
      RECT  139.02 0.62 140.84 1.66 ;
      RECT  142.42 0.62 142.88 1.66 ;
      RECT  151.26 0.62 153.08 1.66 ;
      RECT  154.66 0.62 155.8 1.66 ;
      RECT  168.94 0.62 172.12 1.66 ;
      RECT  181.18 0.62 184.36 1.66 ;
      RECT  191.38 0.62 191.84 1.66 ;
      RECT  193.42 0.62 196.6 1.66 ;
      RECT  204.3 0.62 204.76 1.66 ;
      RECT  206.34 0.62 208.16 1.66 ;
      RECT  215.18 0.62 217.0 1.66 ;
      RECT  218.58 0.62 219.04 1.66 ;
      RECT  227.42 0.62 229.24 1.66 ;
      RECT  230.82 0.62 231.28 1.66 ;
      RECT  238.98 0.62 240.8 1.66 ;
      RECT  242.38 0.62 242.84 1.66 ;
      RECT  249.86 0.62 254.4 1.66 ;
      RECT  268.9 0.62 271.4 1.66 ;
      RECT  281.14 0.62 284.32 1.66 ;
      RECT  291.34 0.62 291.8 1.66 ;
      RECT  293.38 0.62 295.2 1.66 ;
      RECT  296.78 0.62 304.04 1.66 ;
      RECT  305.62 0.62 316.96 1.66 ;
      RECT  318.54 0.62 329.2 1.66 ;
      RECT  330.78 0.62 340.76 1.66 ;
      RECT  342.34 0.62 354.36 1.66 ;
      RECT  355.94 0.62 366.6 1.66 ;
      RECT  368.18 0.62 378.84 1.66 ;
      RECT  380.42 0.62 391.76 1.66 ;
      RECT  393.34 0.62 404.0 1.66 ;
      RECT  405.58 0.62 416.92 1.66 ;
      RECT  418.5 0.62 429.16 1.66 ;
      RECT  430.74 0.62 442.08 1.66 ;
      RECT  443.66 0.62 454.32 1.66 ;
      RECT  455.9 0.62 466.56 1.66 ;
      RECT  468.14 0.62 478.8 1.66 ;
      RECT  480.38 0.62 491.72 1.66 ;
      RECT  493.3 0.62 503.96 1.66 ;
      RECT  505.54 0.62 516.2 1.66 ;
      RECT  517.78 0.62 529.12 1.66 ;
      RECT  530.7 0.62 615.48 1.66 ;
      RECT  116.58 414.88 142.88 415.92 ;
      RECT  144.46 414.88 154.44 415.92 ;
      RECT  156.02 414.88 166.68 415.92 ;
      RECT  168.26 414.88 180.28 415.92 ;
      RECT  181.86 414.88 191.84 415.92 ;
      RECT  193.42 414.88 204.76 415.92 ;
      RECT  206.34 414.88 217.0 415.92 ;
      RECT  218.58 414.88 229.92 415.92 ;
      RECT  231.5 414.88 242.16 415.92 ;
      RECT  243.74 414.88 255.08 415.92 ;
      RECT  256.66 414.88 267.32 415.92 ;
      RECT  268.9 414.88 280.24 415.92 ;
      RECT  281.82 414.88 291.8 415.92 ;
      RECT  293.38 414.88 304.04 415.92 ;
      RECT  305.62 414.88 317.64 415.92 ;
      RECT  319.22 414.88 329.88 415.92 ;
      RECT  331.46 414.88 342.12 415.92 ;
      RECT  343.7 414.88 354.36 415.92 ;
      RECT  355.94 414.88 367.28 415.92 ;
      RECT  368.86 414.88 378.84 415.92 ;
      RECT  380.42 414.88 392.44 415.92 ;
      RECT  394.02 414.88 404.68 415.92 ;
      RECT  406.26 414.88 416.92 415.92 ;
      RECT  418.5 414.88 429.16 415.92 ;
      RECT  430.74 414.88 441.4 415.92 ;
      RECT  442.98 414.88 454.32 415.92 ;
      RECT  455.9 414.88 467.24 415.92 ;
      RECT  468.82 414.88 479.48 415.92 ;
      RECT  481.06 414.88 491.72 415.92 ;
      RECT  493.3 414.88 504.64 415.92 ;
      RECT  506.22 414.88 516.2 415.92 ;
      RECT  517.78 414.88 529.8 415.92 ;
      RECT  531.38 414.88 591.68 415.92 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 412.38 7.1 415.92 ;
      RECT  7.1 1.66 115.0 4.16 ;
      RECT  7.1 4.16 115.0 412.38 ;
      RECT  7.1 412.38 115.0 415.92 ;
      RECT  599.38 1.66 676.0 4.16 ;
      RECT  599.38 4.16 676.0 412.38 ;
      RECT  599.38 412.38 676.0 414.88 ;
      RECT  676.0 1.66 678.94 4.16 ;
      RECT  676.0 412.38 678.94 414.88 ;
      RECT  617.74 0.62 679.4 0.76 ;
      RECT  617.74 0.76 679.4 1.66 ;
      RECT  679.4 0.62 682.34 0.76 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 1.66 ;
      RECT  655.14 414.88 679.4 415.78 ;
      RECT  655.14 415.78 679.4 415.92 ;
      RECT  679.4 415.78 682.34 415.92 ;
      RECT  682.34 414.88 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  678.94 1.66 679.4 4.16 ;
      RECT  682.34 1.66 682.48 4.16 ;
      RECT  678.94 4.16 679.4 412.38 ;
      RECT  682.34 4.16 682.48 412.38 ;
      RECT  678.94 412.38 679.4 414.88 ;
      RECT  682.34 412.38 682.48 414.88 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 79.64 0.76 ;
      RECT  3.7 0.76 79.64 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 412.38 ;
      RECT  3.7 4.16 4.16 412.38 ;
      RECT  0.62 412.38 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 415.78 3.7 415.92 ;
      RECT  3.7 412.38 4.16 415.78 ;
      RECT  3.7 415.78 4.16 415.92 ;
   END
END    sky130_sram_2kbyte_1rw1r_32x512_8
END    LIBRARY
